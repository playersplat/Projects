module countones
  #(parameter width_p = 8)
  (input [width_p - 1:0] binary_i
  ,output [$clog2(width_p) :0] count_o);

  logic [$clog2(width_p) :0] count_l; 

  // For extra credit (25% of Lab 3/Part 3): 
  // 
  // Re-write this loop to synthesize into better hardware. You may
  // not use the $countones() function (though it is synthesizable).
  // 
  // Demonstrate your improvement using the Yosys commands in Piazza.
  always_comb begin
     count_l = 0;
     for(logic [31:0] i = 0; i < width_p; i++) begin
        count_l += {{$clog2(width_p-1){1'b0}},binary_i[i]};
     end
  end
  assign count_o = count_l;

  // Write your immediate and concurrent assertions here

  // The synthesized code below does not implement the correct
  // behavior (but the error is simple).
  // 
  // You must write two concurrent assertions, one demonstrating your understanding
  //
  //  - One must fail (Demonstrating your understanding of how to
  //  write a concurrent assertion that checks for correct behavior.)
  //
  //  - One must pass (Demonstrating your understanding of the bug)
  //

  // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL
 assert property (count_o == $countones(binary_i));
 assert property (count_o == ($countones(binary_i) & {1'bx, 4'b0}));
`endif

endmodule


module countones_synth
  #(parameter width_p = 8)
  (input [width_p - 1:0] binary_i
  ,output [$clog2(width_p) :0] count_o);

  // Write your immediate and concurrent assertions here

  // The synthesized code below does not implement the correct
  // behavior (but the error is simple).
  // 
  // You must write two concurrent assertions, one demonstrating your understanding
  //
  //  - One must fail (Demonstrating your understanding of how to
  //  write a concurrent assertion that checks for correct behavior.)
  //
  //  - One must pass (Demonstrating your understanding of the bug)
  //

  // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL
 assert property (count_o == $countones(binary_i));
 assert property (count_o == ($countones(binary_i) & {1'bx, 4'b0}));
`endif

  yosys_countones
    #()
  countones_synth_i
    (.binary_i(binary_i)
    ,.count_o(count_o));

endmodule


/* Generated by Yosys 0.25 (git sha1 e02b7f64bc7, clang 14.0.0 -fPIC -Os) */

(* hdlname = "\\countones" *)
(* dynports =  1  *)
(* top =  1  *)
(* src = "countones.sv:1.1-40.10" *)
module yosys_countones(binary_i, count_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  (* src = "countones.sv:3.26-3.34" *)
  input [7:0] binary_i;
  wire [7:0] binary_i;
  (* src = "countones.sv:6.30-6.37" *)
  wire [3:0] count_l;
  (* src = "countones.sv:4.32-4.39" *)
  output [3:0] count_o;
  wire [3:0] count_o;
  assign _00_ = ~(binary_i[1] | binary_i[0]);
  assign _01_ = ~binary_i[3];
  assign _02_ = ~(binary_i[1] ^ binary_i[0]);
  assign _03_ = _01_ & ~(_02_);
  assign _04_ = _03_ | _00_;
  assign _05_ = _02_ ^ _01_;
  assign _06_ = _05_ | binary_i[6];
  assign _07_ = ~binary_i[5];
  assign _08_ = ~(_05_ ^ binary_i[6]);
  assign _09_ = _07_ & ~(_08_);
  assign _10_ = _06_ & ~(_09_);
  assign _11_ = _10_ ^ _04_;
  assign _12_ = _08_ ^ _07_;
  assign _13_ = _12_ | binary_i[4];
  assign _14_ = ~binary_i[7];
  assign _15_ = ~(_12_ ^ binary_i[4]);
  assign _16_ = _14_ & ~(_15_);
  assign _17_ = _13_ & ~(_16_);
  assign _18_ = _17_ ^ _11_;
  assign _19_ = _15_ ^ _14_;
  assign _20_ = _19_ | binary_i[2];
  assign count_o[1] = ~(_20_ ^ _18_);
  assign _21_ = _04_ & ~(_10_);
  assign _22_ = _17_ | _11_;
  assign _23_ = _18_ & ~(_20_);
  assign _24_ = _22_ & ~(_23_);
  assign count_o[2] = ~(_24_ ^ _21_);
  assign count_o[0] = _19_ ^ binary_i[2];
  assign count_o[3] = _21_ & ~(_24_);
  assign count_l = count_o;
endmodule

module divider
  #(parameter width_p = 4)
  (input [width_p - 1:0] a_i
  ,input [width_p - 1:0] b_i
  ,output [width_p - 1:0] quot_o
  ,output [width_p - 1:0] rem_o);

  assign quot_o = a_i / b_i;
  assign rem_o = a_i % b_i;

  // Write your immediate and concurrent assertions here

  // The synthesized code below does not implement the correct
  // behavior (but the error is simple).
  // 
  // You must write two concurrent assertions, one demonstrating your understanding
  //
  //  - One must fail (Demonstrating your understanding of how to
  //  write a concurrent assertion that checks for correct behavior.)
  //
  //  - One must pass (Demonstrating your understanding of the bug)
  //

  // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL
 assert property ((quot_o == a_i / b_i) && (rem_o == a_i % b_i));
 assert property (quot_o == ((a_i / b_i) && (rem_o != a_i / b_i))); //test to see if quot_o and rem_o have their logic swapped
`endif

endmodule

module divider_synth
  #(parameter width_p = 4)
  (input [width_p - 1:0] a_i
  ,input [width_p - 1:0] b_i
  ,output [width_p - 1:0] quot_o
  ,output [width_p - 1:0] rem_o);

  // Write your immediate and concurrent assertions here

  // The synthesized code below does not implement the correct
  // behavior (but the error is simple).
  // 
  // You must write two concurrent assertions, one demonstrating your understanding
  //
  //  - One must fail (Demonstrating your understanding of how to
  //  write a concurrent assertion that checks for correct behavior.)
  //
  //  - One must pass (Demonstrating your understanding of the bug)
  //

  // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL
 assert property ((quot_o == a_i / b_i) && (rem_o == a_i % b_i));
 assert property (quot_o == ((a_i / b_i) && (rem_o != a_i / b_i))); //test to see if quot_o and rem_o have their logic swapped
`endif

  yosys_divider
    #()
  divider_synth_i
    (.a_i(a_i)
    ,.b_i(b_i)
    ,.quot_o(quot_o)
    ,.rem_o(rem_o));

endmodule

/* Generated by Yosys 0.25 (git sha1 e02b7f64bc7, clang 14.0.0 -fPIC -Os) */

(* hdlname = "\\divider" *)
(* dynports =  1  *)
(* top =  1  *)
(* src = "divider.sv:1.1-29.10" *)
module yosys_divider(a_i, b_i, quot_o, rem_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  (* src = "divider.sv:3.26-3.29" *)
  input [3:0] a_i;
  wire [3:0] a_i;
  (* src = "divider.sv:4.26-4.29" *)
  input [3:0] b_i;
  wire [3:0] b_i;
  (* src = "divider.sv:5.27-5.33" *)
  output [3:0] quot_o;
  wire [3:0] quot_o;
  (* src = "divider.sv:6.27-6.32" *)
  output [3:0] rem_o;
  wire [3:0] rem_o;
  assign _009_ = ~a_i[3];
  assign _010_ = b_i[0] ^ a_i[3];
  assign _011_ = ~_010_;
  assign _012_ = _010_ | a_i[2];
  assign _013_ = a_i[1] | a_i[0];
  assign _014_ = _013_ | _012_;
  assign _015_ = b_i[1] | b_i[2];
  assign _016_ = _015_ | b_i[3];
  assign _017_ = _016_ | _014_;
  assign _018_ = ~b_i[3];
  assign _019_ = a_i[3] & ~(b_i[0]);
  assign _020_ = a_i[2] & ~(_010_);
  assign _021_ = _020_ | _019_;
  assign _022_ = _012_ & ~(_021_);
  assign _023_ = _022_ | _015_;
  assign _024_ = _018_ & ~(_023_);
  assign _025_ = _017_ & ~(_024_);
  assign _026_ = _025_ ? _009_ : _011_;
  assign _027_ = ~(b_i[2] | b_i[3]);
  assign _028_ = _026_ ^ b_i[1];
  assign _029_ = b_i[0] ^ a_i[2];
  assign _030_ = ~_029_;
  assign _031_ = ~(_030_ & _028_);
  assign _032_ = _031_ | _013_;
  assign _033_ = _032_ | ~(_027_);
  assign _034_ = ~b_i[1];
  assign _035_ = _034_ & ~(_026_);
  assign _036_ = b_i[0] | ~(a_i[2]);
  assign _037_ = _028_ & ~(_036_);
  assign _038_ = _037_ | _035_;
  assign _039_ = _031_ & ~(_038_);
  assign _040_ = _027_ & ~(_039_);
  assign _041_ = _033_ & ~(_040_);
  assign _042_ = b_i[0] & ~(a_i[2]);
  assign _043_ = _042_ ^ _028_;
  assign _044_ = _041_ ? _026_ : _043_;
  assign _045_ = _044_ ^ b_i[2];
  assign _046_ = ~a_i[2];
  assign _047_ = _041_ ? _046_ : _030_;
  assign _048_ = _047_ ^ _034_;
  assign _049_ = _045_ & ~(_048_);
  assign _050_ = b_i[0] ^ a_i[1];
  assign _051_ = ~(_050_ | a_i[0]);
  assign _052_ = ~(_051_ & _049_);
  assign _053_ = _052_ | b_i[3];
  assign _054_ = _044_ | b_i[2];
  assign _055_ = _047_ | b_i[1];
  assign _056_ = _045_ & ~(_055_);
  assign _057_ = _054_ & ~(_056_);
  assign _058_ = b_i[0] & ~(a_i[1]);
  assign _059_ = _049_ & ~(_058_);
  assign _060_ = _057_ & ~(_059_);
  assign _061_ = _018_ & ~(_060_);
  assign _062_ = _053_ & ~(_061_);
  assign _063_ = ~(_058_ | _048_);
  assign _064_ = _055_ & ~(_063_);
  assign _065_ = _064_ ^ _045_;
  assign _066_ = _062_ ? _044_ : _065_;
  assign _067_ = _066_ ^ b_i[3];
  assign _068_ = ~(_058_ ^ _048_);
  assign _069_ = _062_ ? _047_ : _068_;
  assign _070_ = ~(_069_ ^ b_i[2]);
  assign _071_ = _067_ & ~(_070_);
  assign _072_ = ~a_i[1];
  assign _073_ = ~_050_;
  assign _074_ = _062_ ? _072_ : _073_;
  assign _075_ = _074_ ^ _034_;
  assign _076_ = b_i[0] ^ a_i[0];
  assign _077_ = _076_ | _075_;
  assign _078_ = _077_ | ~(_071_);
  assign _079_ = _018_ & ~(_066_);
  assign _080_ = _069_ | b_i[2];
  assign _081_ = _067_ & ~(_080_);
  assign _082_ = _081_ | _079_;
  assign _083_ = _074_ | b_i[1];
  assign _084_ = b_i[0] & ~(a_i[0]);
  assign _085_ = ~(_084_ | _075_);
  assign _086_ = _083_ & ~(_085_);
  assign _087_ = _071_ & ~(_086_);
  assign _088_ = _087_ | _082_;
  assign rem_o[0] = _088_ | ~(_078_);
  assign rem_o[1] = ~_062_;
  assign rem_o[2] = ~_041_;
  assign rem_o[3] = ~_025_;
  assign _000_ = ~_074_;
  assign _001_ = _078_ & ~(_088_);
  assign _002_ = _084_ ^ _075_;
  assign quot_o[1] = _001_ ? _000_ : _002_;
  assign _003_ = ~_069_;
  assign _004_ = _086_ ^ _070_;
  assign quot_o[2] = _001_ ? _003_ : _004_;
  assign quot_o[0] = _001_ ? a_i[0] : _076_;
  assign _005_ = ~_066_;
  assign _006_ = ~(_086_ | _070_);
  assign _007_ = _006_ | ~(_080_);
  assign _008_ = _007_ ^ _067_;
  assign quot_o[3] = _001_ ? _005_ : _008_;
endmodule
